/*
  Yiheng Chi
  chi14@purdue.edu

  hazard control unit test bench
*/

// interface
`include "hazard_control_unit_if.vh"
