/*
  Yiheng Chi
  chi14@purdue.edu

  control unit test bench
*/

// interface
`include "control_unit_if.vh"

// types
`include "cpu_types_pkg.vh"
`include "control_unit_types_pkg.vh"

// mapped timing needs this
`timescale 1 ns / 1 ns

module control_unit_tb;

  // clock period
  parameter PERIOD = 10;

endmodule


