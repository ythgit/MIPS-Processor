/*
  Yiheng Chi
  chi14@purdue.edu

  control unit source code
*/

//
